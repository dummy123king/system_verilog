class  Base;
    int k;
    virtual function void print();
        
    endfunction //new()
endclass // Base


class Derived extends Base;
    virtual function void print();
        
    endfunction //new()
endclass //Derived 